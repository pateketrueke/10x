# Definitions

Local functions can be achieved too:

sum(a, b)=a + b;
sum(1, 2)
