# Maths

Basic operators wors as expected: 1 + 2

Consecutive numbers are always operated, e.g. 1 2 3

# Precedence

Parentheses after numbers are multiplied: 1.5 (2.5 3.5)

The last used operator, plus or minus, is used: 1 2 / 3 - 4 5

You can group expressions within parentheses, e.g. 1 + (2 + 3) / 4 5

# Usage with lists

Same rules applies for numbers inside parentheses and lists, e.g. (1 2 3)

Lists can be mixed, as they aways evaluate expressions inside:

a) (1, 2, 3), 3/2
b) 1 2 / 3, 4 * 5 / 1.5 as fr
c) (1 2) / 3.33 as fr, 4 * 5 / 3 2 as fr
